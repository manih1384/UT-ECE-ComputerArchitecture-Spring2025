module Plus1 (
    input wire [4:0] pc,
    output [4:0] out        
);

assign out = pc+1;

endmodule
