module Plus4 (
    input wire [4:0] pc,
    output [4:0] out        
);

assign out = pc+4;

endmodule
